`ifndef MY_IF__SV
`define MY_IF__SV

interface my_if();
logic[2:0] addr;
data dad;

function void fun1();

endfunction


task dog();

endtask


modport mod1();


clocking clkb@();

endclocking


endinterface
`endif
